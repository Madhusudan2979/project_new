`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 20.10.2023 12:19:39
// Design Name: 
// Module Name: PRNG
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////////////////////////////////////////////////////////////////
module PRNG (
  input logic A,
  input logic clk,
    output logic [11:0] y
);
  logic [11:0]counter1;
  logic [11:0]counter2;
  logic [11:0]a,b,x;
  assign x=8'b11101000;
 initial y=12'b000000000000; 
logic [27:0] counter;
always@(posedge clk)
if (counter[27]==1)
begin 
 counter<=0;
 end 
else
begin 
 counter<=counter+1; 
 end
always_ff @(posedge counter[27]) begin
    if (counter1 < 2047)
      counter1 <= counter1 + 1;
    else
      counter1 <= 0;
  end

  always_ff @(posedge counter[27]) begin
    if (counter2 < 999)
      counter2 <= counter2 + 1;
    else
      counter2 <= 0;
  end

  always_ff@(a, b)
  begin
    a <= counter1[11:0];
    b <= counter2[11:0];
    y <= (a*x+b)%1024;
    end 
endmodule























































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































